module app

import maps
import time
