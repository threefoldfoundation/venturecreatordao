module app

import time

interface IActivity {
	created_at time.Time
}
