module webui
